

module alu (
output reg [31:0] alu_out,
output z,
output reg c,
input [2:0] opcode,
input [31:0] op1,
input [31:0] op2,
input sub
);
reg [31:0] slt_data,sltu_data,srl_data; 

reg [31:0] reg1,reg2;





assign z=~(|alu_out);
parameter 	ADD1 =3'b000,
				SLL1 =3'b001,
				SLT1 =3'b010,
				SLTU1 =3'b011,
				XOR1 =3'b100,
				SRL1 =3'b101,
				OR1 =3'b110,
				AND1 =3'b111;

always@(*)
case(opcode)
		3'b000: {c,alu_out}=(sub==0)?op1+op2:op1-op2;
		3'b110: alu_out=op1|op2;
		3'b100: alu_out=op1^op2;
		3'b111: alu_out=op1&op2;
		3'b001: alu_out=op1<<op2[4:0];
		3'b101: alu_out=srl_data;
		3'b010: alu_out=slt_data;
		3'b011: alu_out=sltu_data;
		default: alu_out={32{1'bx}};
endcase

always@(*)
	if(sub==0)
	srl_data=op1>>op2[4:0];
	else
		begin
			if(op1[31]==1)
				begin
					srl_data=reg1|reg2;
				end
			else
				srl_data=op1>>op2[4:0];
		end
		
always@(*)
	if(op2 > op1)
		sltu_data={{31{1'b0}},1'b1};
	else
		sltu_data=0;
		
always@(*)
	if(op2[31]==1 && op1[31]==0)
		slt_data=0;
	else if(op2[31]==0 && op1[31]==1)
		slt_data={{31{1'b0}},1'b1};
	else if(op2[31]==0 && op1[31]==0)
		begin
				if(op2 > op1)
					slt_data={{31{1'b0}},1'b1};
				else
					slt_data=0;
		end
	else 
		begin
			if(op2[30:0] > op1[30:0])
					slt_data={{31{1'b0}},1'b1};
			else
					slt_data=0;
		end

always@(*)
    case(op2[4:0])    
    5'b00000 :reg1=32'b10000000000000000000000000000000;
    5'b00001 :reg1=32'b11000000000000000000000000000000;
    5'b00010 :reg1=32'b11100000000000000000000000000000;
    5'b00011 :reg1=32'b11110000000000000000000000000000;
    5'b00100 :reg1=32'b11111000000000000000000000000000;
    5'b00101 :reg1=32'b11111100000000000000000000000000;
    5'b00110 :reg1=32'b11111110000000000000000000000000;
    5'b00111 :reg1=32'b11111111000000000000000000000000;
    5'b01000 :reg1=32'b11111111100000000000000000000000;
    5'b01001 :reg1=32'b11111111110000000000000000000000;
    5'b01010 :reg1=32'b11111111111000000000000000000000;
    5'b01011 :reg1=32'b11111111111100000000000000000000;
    5'b01100 :reg1=32'b11111111111110000000000000000000;
    5'b01101 :reg1=32'b11111111111111000000000000000000;
    5'b01110 :reg1=32'b11111111111111100000000000000000;
    5'b01111 :reg1=32'b11111111111111110000000000000000;
    5'b10000 :reg1=32'b11111111111111111000000000000000;
    5'b10001 :reg1=32'b11111111111111111100000000000000;
    5'b10010 :reg1=32'b11111111111111111110000000000000;
    5'b10011 :reg1=32'b11111111111111111111000000000000;
    5'b10100 :reg1=32'b11111111111111111111100000000000;
    5'b10101 :reg1=32'b11111111111111111111110000000000;
    5'b10110 :reg1=32'b11111111111111111111111000000000;
    5'b10111 :reg1=32'b11111111111111111111111100000000;
    5'b11000 :reg1=32'b11111111111111111111111110000000;
    5'b11001 :reg1=32'b11111111111111111111111111000000;
    5'b11010 :reg1=32'b11111111111111111111111111100000;
    5'b11011 :reg1=32'b11111111111111111111111111110000;
    5'b11100 :reg1=32'b11111111111111111111111111111000;
    5'b11101 :reg1=32'b11111111111111111111111111111100;
    5'b11110 :reg1=32'b11111111111111111111111111111110;
    5'b11111 :reg1=32'b11111111111111111111111111111111;
	 default: reg1={32{1'bx}};
endcase

always@(*)
    reg2=op1>>op2[4:0];
    
endmodule  

